/* test for half adder.v 
saved in file half_adder_tb.v*/
`include "half_adder.v"

module half_adder_tb;
 reg a , b; // reg mean register.
 wire sum, carry;
 
 half_adder add1(a,b,sum,carry);

/* code in the initial block executed once
in the entire simulation . Since we have small circuit. it is enough.
begin and end is needed for more than one line of statement.
*/
 initial 
 begin
    $dumpfile("half_adder.vcd"); // value change dump.
    $dumpvars(0,half_adder_tb); 

     a= 0; b = 0;
     #1
     a = 0;b = 1;
     #1
     a = 1;b = 0;
     #1
     a = 1;b = 1;
      
 end
endmodule